
`ifndef ISSUELS_V
`define ISSIELS_V

module issuels (
   input             clk,
   input             reset
);

endmodule

`endif

