
`ifndef IDECODER_V
`define IDECODER_V

module idecoder();


endmodule

`endif

