
`ifndef DIVIDER_V
`define DIVIDER_V

module divider();
endmodule

`endif

