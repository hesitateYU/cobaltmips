-------------------------------------------------------------------------------
--
-- Design       : sprom 
-- Project      : Digilent Terminal 
-- Author       : Srinivas Vaduvatha 
-- Company      : University of Southern California 
--
-------------------------------------------------------------------------------
--
-- File         : sprom.vhd
-- Version      : 1.0
--
-------------------------------------------------------------------------------
--
-- Description  : Data width & Address width - Generics
--                Single port synchronous memory. 
--                Infers BRAM resource in Xilinx FPGAs.
--                If the width / depth specified require more bits than in a single 
--                BRAM, multiple BRAMs are automatically cascaded to form a larger 
--                memory. Memory has to be of (2**n) depth
--
-------------------------------------------------------------------------------

-- libraries and use clauses
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity instruction_mem is 
generic (
         DATA_WIDTH     : integer := 32; 
         ADDR_WIDTH     : integer := 8
        );
port (
      clk           : in  std_logic; 
		en		 		  : in  std_logic;
      addr          : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
      data_out      : out std_logic_vector(DATA_WIDTH-1 downto 0)
     ); 
end instruction_mem ; 

architecture inferrable of instruction_mem is 

-- type declarations
type mem_type is array (0 to(2**ADDR_WIDTH)-1) of std_logic_vector((DATA_WIDTH-1) downto 0); 

-- signals declarations.
signal mem          : mem_type := (X"00422825",X"8C040010",X"00A52820",X"1085fffe",X"00842020",X"00A42024",X"00000020",X"10040004",X"00443020",X"8C030040",X"00642024",X"00642024",X"10C3FFF8",X"00C23022",X"10C5FFFE",X"8CC60010",
											  X"8CC60010",X"10C3FFFC",X"AFA20046",X"00421020",X"00421020",X"00422020",X"00820820",X"AFA1003E",X"8FA3003E",X"AFA30042",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",
											  X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"00000020",X"080000FF");
											  

begin 
mem_read: process (clk) 
begin 
    if (clk = '1' and clk'event) then
		if(en = '1') then
        data_out          <= mem(CONV_INTEGER(addr)); 
		end if;
    end if;
end process; 

end inferrable ;
