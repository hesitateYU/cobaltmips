
`ifndef MULTIPLIER_WRAPPER_V
`define MULTIPLIER_WRAPPER_V

module multiplier_wrapper();
endmodule

`endif

